/**
 * Lookup for a pixel for a number.
 */
module number(
	output reg out,
	input wire[1:0] xpos,
	input wire[2:0] ypos,
	input wire[3:0] value,
	input wire clk
);
	always@(posedge clk) begin
case({value, ypos, xpos})
  9'b000000000: out = 1;
  9'b000000001: out = 1;
  9'b000000010: out = 1;
  9'b000000100: out = 1;
  9'b000000101: out = 0;
  9'b000000110: out = 1;
  9'b000001000: out = 1;
  9'b000001001: out = 0;
  9'b000001010: out = 1;
  9'b000001100: out = 1;
  9'b000001101: out = 0;
  9'b000001110: out = 1;
  9'b000010000: out = 1;
  9'b000010001: out = 1;
  9'b000010010: out = 1;
  9'b000100000: out = 0;
  9'b000100001: out = 1;
  9'b000100010: out = 0;
  9'b000100100: out = 1;
  9'b000100101: out = 1;
  9'b000100110: out = 0;
  9'b000101000: out = 0;
  9'b000101001: out = 1;
  9'b000101010: out = 0;
  9'b000101100: out = 0;
  9'b000101101: out = 1;
  9'b000101110: out = 0;
  9'b000110000: out = 0;
  9'b000110001: out = 1;
  9'b000110010: out = 0;
  9'b001000000: out = 1;
  9'b001000001: out = 1;
  9'b001000010: out = 1;
  9'b001000100: out = 0;
  9'b001000101: out = 0;
  9'b001000110: out = 1;
  9'b001001000: out = 1;
  9'b001001001: out = 1;
  9'b001001010: out = 1;
  9'b001001100: out = 1;
  9'b001001101: out = 0;
  9'b001001110: out = 0;
  9'b001010000: out = 1;
  9'b001010001: out = 1;
  9'b001010010: out = 1;
  9'b001100000: out = 1;
  9'b001100001: out = 1;
  9'b001100010: out = 1;
  9'b001100100: out = 0;
  9'b001100101: out = 0;
  9'b001100110: out = 1;
  9'b001101000: out = 1;
  9'b001101001: out = 1;
  9'b001101010: out = 1;
  9'b001101100: out = 0;
  9'b001101101: out = 0;
  9'b001101110: out = 1;
  9'b001110000: out = 1;
  9'b001110001: out = 1;
  9'b001110010: out = 1;
  9'b010000000: out = 1;
  9'b010000001: out = 0;
  9'b010000010: out = 0;
  9'b010000100: out = 1;
  9'b010000101: out = 0;
  9'b010000110: out = 1;
  9'b010001000: out = 1;
  9'b010001001: out = 1;
  9'b010001010: out = 1;
  9'b010001100: out = 0;
  9'b010001101: out = 0;
  9'b010001110: out = 1;
  9'b010010000: out = 0;
  9'b010010001: out = 0;
  9'b010010010: out = 1;
  9'b010100000: out = 1;
  9'b010100001: out = 1;
  9'b010100010: out = 1;
  9'b010100100: out = 1;
  9'b010100101: out = 0;
  9'b010100110: out = 0;
  9'b010101000: out = 1;
  9'b010101001: out = 1;
  9'b010101010: out = 1;
  9'b010101100: out = 0;
  9'b010101101: out = 0;
  9'b010101110: out = 1;
  9'b010110000: out = 1;
  9'b010110001: out = 1;
  9'b010110010: out = 1;
  9'b011000000: out = 1;
  9'b011000001: out = 1;
  9'b011000010: out = 0;
  9'b011000100: out = 1;
  9'b011000101: out = 0;
  9'b011000110: out = 0;
  9'b011001000: out = 1;
  9'b011001001: out = 1;
  9'b011001010: out = 1;
  9'b011001100: out = 1;
  9'b011001101: out = 0;
  9'b011001110: out = 1;
  9'b011010000: out = 1;
  9'b011010001: out = 1;
  9'b011010010: out = 1;
  9'b011100000: out = 1;
  9'b011100001: out = 1;
  9'b011100010: out = 1;
  9'b011100100: out = 0;
  9'b011100101: out = 0;
  9'b011100110: out = 1;
  9'b011101000: out = 0;
  9'b011101001: out = 1;
  9'b011101010: out = 0;
  9'b011101100: out = 0;
  9'b011101101: out = 1;
  9'b011101110: out = 0;
  9'b011110000: out = 0;
  9'b011110001: out = 1;
  9'b011110010: out = 0;
  9'b100000000: out = 1;
  9'b100000001: out = 1;
  9'b100000010: out = 1;
  9'b100000100: out = 1;
  9'b100000101: out = 0;
  9'b100000110: out = 1;
  9'b100001000: out = 1;
  9'b100001001: out = 1;
  9'b100001010: out = 1;
  9'b100001100: out = 1;
  9'b100001101: out = 0;
  9'b100001110: out = 1;
  9'b100010000: out = 1;
  9'b100010001: out = 1;
  9'b100010010: out = 1;
  9'b100100000: out = 1;
  9'b100100001: out = 1;
  9'b100100010: out = 1;
  9'b100100100: out = 1;
  9'b100100101: out = 0;
  9'b100100110: out = 1;
  9'b100101000: out = 1;
  9'b100101001: out = 1;
  9'b100101010: out = 1;
  9'b100101100: out = 0;
  9'b100101101: out = 0;
  9'b100101110: out = 1;
  9'b100110000: out = 0;
  9'b100110001: out = 1;
  9'b100110010: out = 1;
default: out=0;
endcase
	end




endmodule
