
module configloader (
	noe_in);	

	input		noe_in;
endmodule
